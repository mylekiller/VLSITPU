module TPU_functional (
input reset, clk, sync, out_HL,
output ready, error,
input [7:0] input1,
input [7:0] input2,
output [15:0] out
);



endmodule
